module FIFO_TB();

